module labproject(output logic stepsignal,
						output logic stepsignal_2,
						output logic stepsignal_3,
						output logic dir,		//direction for bending
						output logic dir_2,	//direction for cutting
						output logic testsignal,
						output logic [3:0] ct,
						output logic [7:0] leds,
						(* altera_attribute = "-name WEAK_PULL_UP_RESISTOR ON" *)
						output logic [3:0] kpc,
						input logic [3:0] kpr,
						input logic reset_n, FPGA_CLK1_50);
						
	logic clk2kHz ;                  // 2kHz clock for keypad scanning
	logic kphit ;                		// a key is pressed
	logic [3:0] num ;            		// value of pressed key
	logic [31:0] key;			  			// desired length of wire
	logic onOff ;					  		// determines whether button is pressed or not( maybe not needed)
	
	logic delay;
	
	logic [1:0] digit;
	logic [4:0] num_0, num_1, num_2, num_3;
	logic [7:0] leds_0, leds_1, leds_2, leds_3;
	

	
	pll pll0 ( .inclk0(FPGA_CLK1_50), .c0(clk2kHz) ) ;
	
	always_ff @(posedge clk2kHz)
		digit <= digit + 1'b1;
	
	
	//instantiate modules	
	colseq colseq_0 (.kpc, .clk(clk2kHz), .reset_n, .kpr);
	kpdecode kpdecode_0 (.kpc, .kpr, .num, .kphit);
	key2length key2length_0 (.num, .key);
	time_delay time_delay_9 (.delay, .reset_n, .clk(FPGA_CLK1_50), .keyhit(kphit));
	motortest motortest_0 (.num_0, .num_1, .num_2, .num_3, .reset_n, .stepsignal, .stepsignal_2, .stepsignal_3, .key(num), .onOff(kphit), .delay, .clk(FPGA_CLK1_50), .dir, .dir_2);
	decode7 decode7_0 (.increased_num(num_0), .leds(leds_0)); 
	decode7 decode7_1 (.increased_num(num_1), .leds(leds_1)); 
	decode7 decode7_2 (.increased_num(num_2), .leds(leds_2)); 
	decode7 decode7_3 (.increased_num(num_3), .leds(leds_3)); 
	decode2 decode2_0 (.leds, .digit, .ct, .leds_0, .leds_1, .leds_2, .leds_3);

endmodule


// megafunction wizard: %ALTPLL%
// ...
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
// ...

module pll ( inclk0, c0);

        input     inclk0;
        output    c0;

        wire [0:0] sub_wire2 = 1'h0;
        wire [4:0] sub_wire3;
        wire  sub_wire0 = inclk0;
        wire [1:0] sub_wire1 = {sub_wire2, sub_wire0};
        wire [0:0] sub_wire4 = sub_wire3[0:0];
        wire  c0 = sub_wire4;

        altpll altpll_component ( .inclk (sub_wire1), .clk
          (sub_wire3), .activeclock (), .areset (1'b0), .clkbad
          (), .clkena ({6{1'b1}}), .clkloss (), .clkswitch
          (1'b0), .configupdate (1'b0), .enable0 (), .enable1 (),
          .extclk (), .extclkena ({4{1'b1}}), .fbin (1'b1),
          .fbmimicbidir (), .fbout (), .fref (), .icdrclk (),
          .locked (), .pfdena (1'b1), .phasecounterselect
          ({4{1'b1}}), .phasedone (), .phasestep (1'b1),
          .phaseupdown (1'b1), .pllena (1'b1), .scanaclr (1'b0),
          .scanclk (1'b0), .scanclkena (1'b1), .scandata (1'b0),
          .scandataout (), .scandone (), .scanread (1'b0),
          .scanwrite (1'b0), .sclkout0 (), .sclkout1 (),
          .vcooverrange (), .vcounderrange ());

        defparam
                altpll_component.bandwidth_type = "AUTO",
                altpll_component.clk0_divide_by = 25000,
                altpll_component.clk0_duty_cycle = 50,
                altpll_component.clk0_multiply_by = 1,
                altpll_component.clk0_phase_shift = "0",
                altpll_component.compensate_clock = "CLK0",
                altpll_component.inclk0_input_frequency = 20000,
                altpll_component.intended_device_family = "Cyclone IV E",
                altpll_component.lpm_hint = "CBX_MODULE_PREFIX=lab1clk",
                altpll_component.lpm_type = "altpll",
                altpll_component.operation_mode = "NORMAL",
                altpll_component.pll_type = "AUTO",
                altpll_component.port_activeclock = "PORT_UNUSED",
                altpll_component.port_areset = "PORT_UNUSED",
                altpll_component.port_clkbad0 = "PORT_UNUSED",
                altpll_component.port_clkbad1 = "PORT_UNUSED",
                altpll_component.port_clkloss = "PORT_UNUSED",
                altpll_component.port_clkswitch = "PORT_UNUSED",
                altpll_component.port_configupdate = "PORT_UNUSED",
                altpll_component.port_fbin = "PORT_UNUSED",
                altpll_component.port_inclk0 = "PORT_USED",
                altpll_component.port_inclk1 = "PORT_UNUSED",
                altpll_component.port_locked = "PORT_UNUSED",
                altpll_component.port_pfdena = "PORT_UNUSED",
                altpll_component.port_phasecounterselect = "PORT_UNUSED",
                altpll_component.port_phasedone = "PORT_UNUSED",
                altpll_component.port_phasestep = "PORT_UNUSED",
                altpll_component.port_phaseupdown = "PORT_UNUSED",
                altpll_component.port_pllena = "PORT_UNUSED",
                altpll_component.port_scanaclr = "PORT_UNUSED",
                altpll_component.port_scanclk = "PORT_UNUSED",
                altpll_component.port_scanclkena = "PORT_UNUSED",
                altpll_component.port_scandata = "PORT_UNUSED",
                altpll_component.port_scandataout = "PORT_UNUSED",
                altpll_component.port_scandone = "PORT_UNUSED",
                altpll_component.port_scanread = "PORT_UNUSED",
                altpll_component.port_scanwrite = "PORT_UNUSED",
                altpll_component.port_clk0 = "PORT_USED",
                altpll_component.port_clk1 = "PORT_UNUSED",
                altpll_component.port_clk2 = "PORT_UNUSED",
                altpll_component.port_clk3 = "PORT_UNUSED",
                altpll_component.port_clk4 = "PORT_UNUSED",
                altpll_component.port_clk5 = "PORT_UNUSED",
                altpll_component.port_clkena0 = "PORT_UNUSED",
                altpll_component.port_clkena1 = "PORT_UNUSED",
                altpll_component.port_clkena2 = "PORT_UNUSED",
                altpll_component.port_clkena3 = "PORT_UNUSED",
                altpll_component.port_clkena4 = "PORT_UNUSED",
                altpll_component.port_clkena5 = "PORT_UNUSED",
                altpll_component.port_extclk0 = "PORT_UNUSED",
                altpll_component.port_extclk1 = "PORT_UNUSED",
                altpll_component.port_extclk2 = "PORT_UNUSED",
                altpll_component.port_extclk3 = "PORT_UNUSED",
                altpll_component.width_clock = 5;


endmodule
