module labproject(output logic [35:0] GPIO_1);
	
	assign GPIO_1[0] = 1'b1;

endmodule